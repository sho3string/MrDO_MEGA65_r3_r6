----------------------------------------------------------------------------------
-- MiSTer2MEGA65 Framework
--
-- Global constants
--
-- MiSTer2MEGA65 done by sy2002 and MJoergen in 2022 and licensed under GPL v3
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.NUMERIC_STD_UNSIGNED.ALL;

library work;
use work.qnice_tools.all;
use work.video_modes_pkg.all;

package globals is

----------------------------------------------------------------------------------------------------------
-- QNICE Firmware
----------------------------------------------------------------------------------------------------------

-- QNICE Firmware: Use the regular QNICE "operating system" called "Monitor" while developing and
-- debugging the firmware/ROM itself. If you are using the M2M ROM (the "Shell") as provided by the
-- framework, then always use the release version of the M2M firmware: QNICE_FIRMWARE_M2M
--
-- Hint: You need to run QNICE/tools/make-toolchain.sh to obtain "monitor.rom" and
-- you need to run CORE/m2m-rom/make_rom.sh to obtain the .rom file
constant QNICE_FIRMWARE_MONITOR   : string  := "../../../M2M/QNICE/monitor/monitor.rom";    -- debug/development
constant QNICE_FIRMWARE_M2M       : string  := "../../../CORE/m2m-rom/m2m-rom.rom";         -- release

-- Select firmware here
constant QNICE_FIRMWARE           : string  := QNICE_FIRMWARE_M2M;

----------------------------------------------------------------------------------------------------------
-- Clock Speed(s)
--
-- Important: Make sure that you use very exact numbers - down to the actual Hertz - because some cores
-- rely on these exact numbers. By default M2M supports one core clock speed. In case you need more,
-- then add all the clocks speeds here by adding more constants.
----------------------------------------------------------------------------------------------------------

-- Galaga core's clock speed
-- Actual clock is 49 Mhz ( see MAME driver - MrDo.cpp ).
-- MiSTer uses 18Mhz
constant CORE_CLK_SPEED       : natural := 49_000_000;   -- Mr Do's main & video clock is 49 MHz 

-- System clock speed (crystal that is driving the FPGA) and QNICE clock speed
-- !!! Do not touch !!!
constant BOARD_CLK_SPEED      : natural := 100_000_000;
constant QNICE_CLK_SPEED      : natural := 50_000_000;   -- a change here has dependencies in qnice_globals.vhd

----------------------------------------------------------------------------------------------------------
-- Video Mode
----------------------------------------------------------------------------------------------------------

-- Rendering constants (in pixels)
--    VGA_*   size of the core's target output post scandoubler
--    FONT_*  size of one OSM character
constant VGA_DX               : natural := 496;
constant VGA_DY               : natural := 384;
constant FONT_FILE            : string  := "../font/Anikki-16x16-m2m.rom";
constant FONT_DX              : natural := 16;
constant FONT_DY              : natural := 16;

-- Constants for the OSM screen memory
constant CHARS_DX             : natural := VGA_DX / FONT_DX;
constant CHARS_DY             : natural := VGA_DY / FONT_DY;
constant CHAR_MEM_SIZE        : natural := CHARS_DX * CHARS_DY;
constant VRAM_ADDR_WIDTH      : natural := f_log2(CHAR_MEM_SIZE);

----------------------------------------------------------------------------------------------------------
-- HyperRAM memory map (in units of 4kW)
----------------------------------------------------------------------------------------------------------

constant C_HMAP_M2M           : std_logic_vector(15 downto 0) := x"0000";     -- Reserved for the M2M framework
constant C_HMAP_DEMO          : std_logic_vector(15 downto 0) := x"0200";     -- Start address reserved for core

----------------------------------------------------------------------------------------------------------
-- Virtual Drive Management System
----------------------------------------------------------------------------------------------------------

-- Virtual drive management system (handled by vdrives.vhd and the firmware)
-- If you are not using virtual drives, make sure that:
--    C_VDNUM        is 0
--    C_VD_DEVICE    is x"EEEE"
--    C_VD_BUFFER    is (x"EEEE", x"EEEE")
-- Otherwise make sure that you wire C_VD_DEVICE in the qnice_ramrom_devices process and that you
-- have as many appropriately sized RAM buffers for disk images as you have drives
type vd_buf_array is array(natural range <>) of std_logic_vector;
constant C_VDNUM              : natural := 0;
constant C_VD_DEVICE          : std_logic_vector(15 downto 0) := x"EEEE";
constant C_VD_BUFFER          : vd_buf_array := (x"EEEE", x"EEEE");

----------------------------------------------------------------------------------------------------------
-- System for handling simulated cartridges and ROM loaders
----------------------------------------------------------------------------------------------------------

type crtrom_buf_array is array(natural range<>) of std_logic_vector;
constant ENDSTR : character := character'val(0);

-- Cartridges and ROMs can be stored into QNICE devices, HyperRAM and SDRAM
constant C_CRTROMTYPE_DEVICE     : std_logic_vector(15 downto 0) := x"0000";
constant C_CRTROMTYPE_HYPERRAM   : std_logic_vector(15 downto 0) := x"0001";
constant C_CRTROMTYPE_SDRAM      : std_logic_vector(15 downto 0) := x"0002";           -- @TODO/RESERVED for future R4 boards

-- Types of automatically loaded ROMs:
-- If a mandatory file is missing, then the core outputs the missing file and goes fatal
constant C_CRTROMTYPE_MANDATORY  : std_logic_vector(15 downto 0) := x"0003";
constant C_CRTROMTYPE_OPTIONAL   : std_logic_vector(15 downto 0) := x"0004";


-- Manually loadable ROMs and cartridges as defined in config.vhd
-- If you are not using this, then make sure that:
--    C_CRTROM_MAN_NUM    is 0
--    C_CRTROMS_MAN       is (x"EEEE", x"EEEE", x"EEEE")
-- Each entry of the array consists of two constants:
--    1) Type of CRT or ROM: Load to a QNICE device, load into HyperRAM, load into SDRAM
--    2) If (1) = QNICE device, then this is the device ID
--       else it is a 4k window in HyperRAM or in SDRAM
-- In case we are loading to a QNICE device, then the control and status register is located at the 4k window 0xFFFF.
-- @TODO: See @TODO for more details about the control and status register
constant C_CRTROMS_MAN_NUM       : natural := 0;                                       -- amount of manually loadable ROMs and carts, if more than 3: also adjust CRTROM_MAN_MAX in M2M/rom/shell_vars.asm, Needs to be in sync with config.vhd. Maximum is 16
constant C_CRTROMS_MAN           : crtrom_buf_array := ( x"EEEE", x"EEEE",
                                                         x"EEEE");                     -- Always finish the array using x"EEEE"

-- Automatically loaded ROMs: These ROMs are loaded before the core starts
--
-- Works similar to manually loadable ROMs and cartridges and each line item has two additional parameters:
--    1) and 2) see above
--    3) Mandatory or optional ROM
--    4) Start address of ROM file name within C_CRTROM_AUTO_NAMES
-- If you are not using this, then make sure that:
--    C_CRTROMS_AUTO_NUM  is 0
--    C_CRTROMS_AUTO      is (x"EEEE", x"EEEE", x"EEEE", x"EEEE", x"EEEE")
-- How to pass the filenames of the ROMs to the framework:
-- C_CRTROMS_AUTO_NAMES is a concatenation of all filenames (see config.vhd's WHS_DATA for an example of how to concatenate)
--    The start addresses of the filename can be determined similarly to how it is done in config.vhd's HELP_x_START
--    using a concatenated addition and VHDL's string length operator.
--    IMPORTANT: a) The framework is not doing any consistency or error check when it comes to C_CRTROMS_AUTO_NAMES, so you
--                  need to be extra careful that the string itself plus the start position of the namex are correct.
--               b) Don't forget to zero-terminate each of your substrings of C_CRTROMS_AUTO_NAMES by adding "& ENDSTR;"
--               c) Don't forget to finish the C_CRTROMS_AUTO array with x"EEEE"

constant C_DEV_A4           : std_logic_vector(15 downto 0) := x"0100"; 
constant C_DEV_C4           : std_logic_vector(15 downto 0) := x"0101";
constant C_DEV_E4           : std_logic_vector(15 downto 0) := x"0102";
constant C_DEV_F4           : std_logic_vector(15 downto 0) := x"0103";
constant C_DEV_S8           : std_logic_vector(15 downto 0) := x"0104";
constant C_DEV_U8           : std_logic_vector(15 downto 0) := x"0105";
constant C_DEV_R8           : std_logic_vector(15 downto 0) := x"0106";
constant C_DEV_N8           : std_logic_vector(15 downto 0) := x"0107";
constant C_DEV_H5           : std_logic_vector(15 downto 0) := x"0108";
constant C_DEV_K5           : std_logic_vector(15 downto 0) := x"0109";
constant C_DEV_U02          : std_logic_vector(15 downto 0) := x"010A";
constant C_DEV_T02          : std_logic_vector(15 downto 0) := x"010B";
constant C_DEV_F10          : std_logic_vector(15 downto 0) := x"010C";


-- Mr Do core specific ROMs
constant ROM_A4             : string  := "arcade/mrdo/a4-01.bin" & ENDSTR;
constant ROM_C4             : string  := "arcade/mrdo/c4-02.bin" & ENDSTR;
constant ROM_E4             : string  := "arcade/mrdo/e4-03.bin" & ENDSTR;
constant ROM_F4             : string  := "arcade/mrdo/f4-04.bin" & ENDSTR;
constant ROM_S8             : string  := "arcade/mrdo/s8-09.bin" & ENDSTR;
constant ROM_U8             : string  := "arcade/mrdo/u8-10.bin" & ENDSTR;
constant ROM_R8             : string  := "arcade/mrdo/r8-08.bin" & ENDSTR;
constant ROM_N8             : string  := "arcade/mrdo/n8-07.bin" & ENDSTR;
constant ROM_H5             : string  := "arcade/mrdo/h5-05.bin" & ENDSTR;
constant ROM_K5             : string  := "arcade/mrdo/k5-06.bin" & ENDSTR;
constant ROM_U02            : string  := "arcade/mrdo/u02--2.bin" & ENDSTR;
constant ROM_T02            : string  := "arcade/mrdo/t02--3.bin" & ENDSTR;
constant ROM_F10            : string  := "arcade/mrdo/f10--1.bin" & ENDSTR;

constant ROM_A4_START          : std_logic_vector(15 downto 0) := X"0000";
constant ROM_C4_START          : std_logic_vector(15 downto 0) := ROM_A4_START + ROM_A4'length;
constant ROM_E4_START          : std_logic_vector(15 downto 0) := ROM_C4_START + ROM_C4'length;
constant ROM_F4_START          : std_logic_vector(15 downto 0) := ROM_E4_START + ROM_E4'length;
constant ROM_S8_START          : std_logic_vector(15 downto 0) := ROM_F4_START + ROM_F4'length;
constant ROM_U8_START          : std_logic_vector(15 downto 0) := ROM_S8_START + ROM_S8'length;
constant ROM_R8_START          : std_logic_vector(15 downto 0) := ROM_U8_START + ROM_U8'length;
constant ROM_N8_START          : std_logic_vector(15 downto 0) := ROM_R8_START + ROM_R8'length;
constant ROM_H5_START          : std_logic_vector(15 downto 0) := ROM_N8_START + ROM_N8'length;
constant ROM_K5_START          : std_logic_vector(15 downto 0) := ROM_H5_START + ROM_H5'length;
constant ROM_U02_START         : std_logic_vector(15 downto 0) := ROM_K5_START + ROM_K5'length;
constant ROM_T02_START         : std_logic_vector(15 downto 0) := ROM_U02_START + ROM_U02'length;
constant ROM_F10_START         : std_logic_vector(15 downto 0) := ROM_T02_START + ROM_T02'length;


-- M2M framework constants
constant C_CRTROMS_AUTO_NUM      : natural := 13;                                       -- Amount of automatically loadable ROMs and carts, if more tha    n 3: also adjust CRTROM_MAN_MAX in M2M/rom/shell_vars.asm, Needs to be in sync with config.vhd. Maximum is 16
constant C_CRTROMS_AUTO_NAMES    : string  := ROM_A4 & ROM_C4 & ROM_E4 & ROM_F4 & 
                                              ROM_S8 & ROM_U8 & ROM_R8 & ROM_N8 &
                                              ROM_H5 & ROM_K5 & ROM_U02 & ROM_T02 & ROM_F10 &
                                              ENDSTR;
                                              
constant C_CRTROMS_AUTO          : crtrom_buf_array := ( 
      C_CRTROMTYPE_DEVICE, C_DEV_A4, C_CRTROMTYPE_MANDATORY, ROM_A4_START,
      C_CRTROMTYPE_DEVICE, C_DEV_C4, C_CRTROMTYPE_MANDATORY, ROM_C4_START,
      C_CRTROMTYPE_DEVICE, C_DEV_E4, C_CRTROMTYPE_MANDATORY, ROM_E4_START,
      C_CRTROMTYPE_DEVICE, C_DEV_F4, C_CRTROMTYPE_MANDATORY, ROM_F4_START,
      C_CRTROMTYPE_DEVICE, C_DEV_S8, C_CRTROMTYPE_MANDATORY, ROM_S8_START,
      C_CRTROMTYPE_DEVICE, C_DEV_U8, C_CRTROMTYPE_MANDATORY, ROM_U8_START,
      C_CRTROMTYPE_DEVICE, C_DEV_R8, C_CRTROMTYPE_MANDATORY, ROM_R8_START,
      C_CRTROMTYPE_DEVICE, C_DEV_N8, C_CRTROMTYPE_MANDATORY, ROM_N8_START,
      C_CRTROMTYPE_DEVICE, C_DEV_H5, C_CRTROMTYPE_MANDATORY, ROM_H5_START,
      C_CRTROMTYPE_DEVICE, C_DEV_K5, C_CRTROMTYPE_MANDATORY, ROM_K5_START,
      C_CRTROMTYPE_DEVICE, C_DEV_U02,C_CRTROMTYPE_MANDATORY, ROM_U02_START,
      C_CRTROMTYPE_DEVICE, C_DEV_T02,C_CRTROMTYPE_MANDATORY, ROM_T02_START,
      C_CRTROMTYPE_DEVICE, C_DEV_F10,C_CRTROMTYPE_MANDATORY, ROM_F10_START,
                                                         x"EEEE");                     -- Always finish the array using x"EEEE"


----------------------------------------------------------------------------------------------------------
-- Audio filters
--
-- If you use audio filters, then you need to copy the correct values from the MiSTer core
-- that you are porting: sys/sys_top.v
----------------------------------------------------------------------------------------------------------

-- Sample values from the C64: @TODO: Adjust to your needs
constant audio_flt_rate : std_logic_vector(31 downto 0) := std_logic_vector(to_signed(7056000, 32));
constant audio_cx       : std_logic_vector(39 downto 0) := std_logic_vector(to_signed(4258969, 40));
constant audio_cx0      : std_logic_vector( 7 downto 0) := std_logic_vector(to_signed(3, 8));
constant audio_cx1      : std_logic_vector( 7 downto 0) := std_logic_vector(to_signed(2, 8));
constant audio_cx2      : std_logic_vector( 7 downto 0) := std_logic_vector(to_signed(1, 8));
constant audio_cy0      : std_logic_vector(23 downto 0) := std_logic_vector(to_signed(-6216759, 24));
constant audio_cy1      : std_logic_vector(23 downto 0) := std_logic_vector(to_signed( 6143386, 24));
constant audio_cy2      : std_logic_vector(23 downto 0) := std_logic_vector(to_signed(-2023767, 24));
constant audio_att      : std_logic_vector( 4 downto 0) := "00000";
constant audio_mix      : std_logic_vector( 1 downto 0) := "00"; -- 0 - no mix, 1 - 25%, 2 - 50%, 3 - 100% (mono)

end package globals;